`define pkt 5
